library ieee;
use ieee.std_logic_1164.all;
entity master is 
    port(
        clk   : in std_logic;     
        reset : in std_logic;     -- Reset signal
        miso  : in std_logic;     -- Master In Slave Out, input from slave
        mosi  : out std_logic;    -- Master Out Slave In, output to slave
        cs    : out std_logic;    -- Chip select, output to slave
        sclk  : out std_logic;
		  data_in : out STD_LOGIC_VECTOR(2 downto 0) := (others => '0')
    );
end entity master;

architecture logic of master is 
    signal sclk_gen : std_logic := '0';    -- SPI clock generated by master
    signal clk_counter   : integer range 0 to 4 := 0;
    signal bit_counter   : integer range 0 to 4 := 0;
    signal datatransmitted : std_logic_vector(2 downto 0) := "101";  -- Data to transmit
    signal cs_gen     : std_logic := '1';  
begin
    -- Clock generation process (SPI clock, SCLK)
    process(clk, reset)
    begin
        if (reset = '1') then
            clk_counter <= 0;
            sclk_gen <= '0';    -- Reset the SPI clock
        elsif rising_edge(clk) then
            if clk_counter = 4 then      -- Divide the system clock by 5
                clk_counter <= 0;
                sclk_gen <= not sclk_gen;  -- Toggle the SPI clock
            else 
                clk_counter <= clk_counter + 1;
            end if;
        end if;
    end process;
	 
    -- Transmitting data (on the falling edge of the SPI clock)
	 
    process(sclk_gen, reset)
    begin
        if reset = '1' then
            mosi <= '0';
            bit_counter <= 0;
				cs_gen <= '1';
        elsif falling_edge(sclk_gen) then  
			   if(bit_counter = 0) then
					cs_gen <= '0';
				end if;
				if(cs_gen = '0') then
					if bit_counter >2 then 
						mosi <= '0';
					end if;
					if(bit_counter < 3) then
						mosi <= datatransmitted(bit_counter);
					end if;
					
					if bit_counter < 4 then
						bit_counter <= bit_counter + 1;
					elsif bit_counter = 4 then
						cs_gen <= '1';
					end if;
				else
						mosi <= '0';
					
            end if;
        end if;
    end process;
	 
	 process(sclk_gen,reset)
	 begin
			if reset ='1' then 
				data_in <= (others => '0');
			elsif rising_edge(SCLK_gen) and bit_counter > 0 then
				if cs_gen = '0' then
					if(bit_counter < 4) then
						data_in(bit_counter-1) <= MISO;
					end if;
				else 
					data_in <= (others => '0');
				end if;
			end if;
	 end process;
    sclk <= sclk_gen;
    cs <= cs_gen;
end architecture logic; 